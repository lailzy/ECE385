module IR(
    input logic Clk,


);
endmodule